// Code your testbench here
// or browse Examples
module fir_filter_pipeline_tb();
reg clk;
reg reset;
reg [15:0] sample;
wire [31:0] result;
wire [31:0] noisy_sample;

fir_filter_pipeline uut(
.clk(clk),
.reset(reset),
.sample(sample),
.result(result),
.noisy_sample(noisy_sample)
);

integer i;
reg [15:0] ecg_samples [0:999]; // array to store ECG samples

initial begin
ecg_samples[0] = 16'd995;
ecg_samples[1] = 16'd995;
ecg_samples[2] = 16'd995;
ecg_samples[3] = 16'd995;
ecg_samples[4] = 16'd995;
ecg_samples[5] = 16'd995;
ecg_samples[6] = 16'd995;
ecg_samples[7] = 16'd995;
ecg_samples[8] = 16'd1000;
ecg_samples[9] = 16'd1000;
ecg_samples[10] = 16'd997;
ecg_samples[11] = 16'd995;
ecg_samples[12] = 16'd994;
ecg_samples[13] = 16'd992;
ecg_samples[14] = 16'd993;
ecg_samples[15] = 16'd992;
ecg_samples[16] = 16'd989;
ecg_samples[17] = 16'd988;
ecg_samples[18] = 16'd987;
ecg_samples[19] = 16'd990;
ecg_samples[20] = 16'd993;
ecg_samples[21] = 16'd989;
ecg_samples[22] = 16'd988;
ecg_samples[23] = 16'd986;
ecg_samples[24] = 16'd988;
ecg_samples[25] = 16'd993;
ecg_samples[26] = 16'd997;
ecg_samples[27] = 16'd993;
ecg_samples[28] = 16'd986;
ecg_samples[29] = 16'd983;
ecg_samples[30] = 16'd977;
ecg_samples[31] = 16'd979;
ecg_samples[32] = 16'd975;
ecg_samples[33] = 16'd974;
ecg_samples[34] = 16'd972;
ecg_samples[35] = 16'd969;
ecg_samples[36] = 16'd969;
ecg_samples[37] = 16'd969;
ecg_samples[38] = 16'd971;
ecg_samples[39] = 16'd973;
ecg_samples[40] = 16'd971;
ecg_samples[41] = 16'd969;
ecg_samples[42] = 16'd966;
ecg_samples[43] = 16'd966;
ecg_samples[44] = 16'd966;
ecg_samples[45] = 16'd966;
ecg_samples[46] = 16'd967;
ecg_samples[47] = 16'd965;
ecg_samples[48] = 16'd963;
ecg_samples[49] = 16'd967;
ecg_samples[50] = 16'd969;
ecg_samples[51] = 16'd969;
ecg_samples[52] = 16'd968;
ecg_samples[53] = 16'd967;
ecg_samples[54] = 16'd963;
ecg_samples[55] = 16'd966;
ecg_samples[56] = 16'd964;
ecg_samples[57] = 16'd968;
ecg_samples[58] = 16'd966;
ecg_samples[59] = 16'd964;
ecg_samples[60] = 16'd961;
ecg_samples[61] = 16'd960;
ecg_samples[62] = 16'd957;
ecg_samples[63] = 16'd952;
ecg_samples[64] = 16'd947;
ecg_samples[65] = 16'd947;
ecg_samples[66] = 16'd943;
ecg_samples[67] = 16'd933;
ecg_samples[68] = 16'd927;
ecg_samples[69] = 16'd927;
ecg_samples[70] = 16'd939;
ecg_samples[71] = 16'd958;
ecg_samples[72] = 16'd980;
ecg_samples[73] = 16'd1010;
ecg_samples[74] = 16'd1048;
ecg_samples[75] = 16'd1099;
ecg_samples[76] = 16'd1148;
ecg_samples[77] = 16'd1180;
ecg_samples[78] = 16'd1192;
ecg_samples[79] = 16'd1177;
ecg_samples[80] = 16'd1128;
ecg_samples[81] = 16'd1058;
ecg_samples[82] = 16'd991;
ecg_samples[83] = 16'd951;
ecg_samples[84] = 16'd937;
ecg_samples[85] = 16'd939;
ecg_samples[86] = 16'd950;
ecg_samples[87] = 16'd958;
ecg_samples[88] = 16'd959;
ecg_samples[89] = 16'd957;
ecg_samples[90] = 16'd955;
ecg_samples[91] = 16'd958;
ecg_samples[92] = 16'd959;
ecg_samples[93] = 16'd961;
ecg_samples[94] = 16'd962;
ecg_samples[95] = 16'd960;
ecg_samples[96] = 16'd957;
ecg_samples[97] = 16'd956;
ecg_samples[98] = 16'd959;
ecg_samples[99] = 16'd955;
ecg_samples[100] = 16'd957;
ecg_samples[101] = 16'd958;
ecg_samples[102] = 16'd957;
ecg_samples[103] = 16'd958;
ecg_samples[104] = 16'd959;
ecg_samples[105] = 16'd958;
ecg_samples[106] = 16'd958;
ecg_samples[107] = 16'd955;
ecg_samples[108] = 16'd953;
ecg_samples[109] = 16'd957;
ecg_samples[110] = 16'd959;
ecg_samples[111] = 16'd963;
ecg_samples[112] = 16'd960;
ecg_samples[113] = 16'd960;
ecg_samples[114] = 16'd958;
ecg_samples[115] = 16'd956;
ecg_samples[116] = 16'd957;
ecg_samples[117] = 16'd956;
ecg_samples[118] = 16'd955;
ecg_samples[119] = 16'd953;
ecg_samples[120] = 16'd953;
ecg_samples[121] = 16'd956;
ecg_samples[122] = 16'd958;
ecg_samples[123] = 16'd958;
ecg_samples[124] = 16'd958;
ecg_samples[125] = 16'd956;
ecg_samples[126] = 16'd954;
ecg_samples[127] = 16'd959;
ecg_samples[128] = 16'd959;
ecg_samples[129] = 16'd958;
ecg_samples[130] = 16'd958;
ecg_samples[131] = 16'd957;
ecg_samples[132] = 16'd957;
ecg_samples[133] = 16'd956;
ecg_samples[134] = 16'd958;
ecg_samples[135] = 16'd956;
ecg_samples[136] = 16'd954;
ecg_samples[137] = 16'd953;
ecg_samples[138] = 16'd954;
ecg_samples[139] = 16'd955;
ecg_samples[140] = 16'd958;
ecg_samples[141] = 16'd960;
ecg_samples[142] = 16'd957;
ecg_samples[143] = 16'd958;
ecg_samples[144] = 16'd955;
ecg_samples[145] = 16'd958;
ecg_samples[146] = 16'd957;
ecg_samples[147] = 16'd957;
ecg_samples[148] = 16'd955;
ecg_samples[149] = 16'd955;
ecg_samples[150] = 16'd953;
ecg_samples[151] = 16'd956;
ecg_samples[152] = 16'd956;
ecg_samples[153] = 16'd957;
ecg_samples[154] = 16'd958;
ecg_samples[155] = 16'd954;
ecg_samples[156] = 16'd954;
ecg_samples[157] = 16'd955;
ecg_samples[158] = 16'd957;
ecg_samples[159] = 16'd957;
ecg_samples[160] = 16'd957;
ecg_samples[161] = 16'd954;
ecg_samples[162] = 16'd953;
ecg_samples[163] = 16'd953;
ecg_samples[164] = 16'd955;
ecg_samples[165] = 16'd955;
ecg_samples[166] = 16'd957;
ecg_samples[167] = 16'd954;
ecg_samples[168] = 16'd952;
ecg_samples[169] = 16'd952;
ecg_samples[170] = 16'd952;
ecg_samples[171] = 16'd951;
ecg_samples[172] = 16'd952;
ecg_samples[173] = 16'd950;
ecg_samples[174] = 16'd947;
ecg_samples[175] = 16'd950;
ecg_samples[176] = 16'd952;
ecg_samples[177] = 16'd953;
ecg_samples[178] = 16'd952;
ecg_samples[179] = 16'd949;
ecg_samples[180] = 16'd949;
ecg_samples[181] = 16'd951;
ecg_samples[182] = 16'd951;
ecg_samples[183] = 16'd952;
ecg_samples[184] = 16'd952;
ecg_samples[185] = 16'd951;
ecg_samples[186] = 16'd950;
ecg_samples[187] = 16'd953;
ecg_samples[188] = 16'd958;
ecg_samples[189] = 16'd959;
ecg_samples[190] = 16'd959;
ecg_samples[191] = 16'd957;
ecg_samples[192] = 16'd956;
ecg_samples[193] = 16'd961;
ecg_samples[194] = 16'd964;
ecg_samples[195] = 16'd964;
ecg_samples[196] = 16'd966;
ecg_samples[197] = 16'd965;
ecg_samples[198] = 16'd966;
ecg_samples[199] = 16'd967;
ecg_samples[200] = 16'd969;
ecg_samples[201] = 16'd973;
ecg_samples[202] = 16'd974;
ecg_samples[203] = 16'd974;
ecg_samples[204] = 16'd971;
ecg_samples[205] = 16'd973;
ecg_samples[206] = 16'd975;
ecg_samples[207] = 16'd978;
ecg_samples[208] = 16'd975;
ecg_samples[209] = 16'd975;
ecg_samples[210] = 16'd973;
ecg_samples[211] = 16'd973;
ecg_samples[212] = 16'd976;
ecg_samples[213] = 16'd974;
ecg_samples[214] = 16'd973;
ecg_samples[215] = 16'd975;
ecg_samples[216] = 16'd973;
ecg_samples[217] = 16'd974;
ecg_samples[218] = 16'd974;
ecg_samples[219] = 16'd971;
ecg_samples[220] = 16'd972;
ecg_samples[221] = 16'd972;
ecg_samples[222] = 16'd971;
ecg_samples[223] = 16'd970;
ecg_samples[224] = 16'd971;
ecg_samples[225] = 16'd972;
ecg_samples[226] = 16'd969;
ecg_samples[227] = 16'd968;
ecg_samples[228] = 16'd966;
ecg_samples[229] = 16'd969;
ecg_samples[230] = 16'd970;
ecg_samples[231] = 16'd972;
ecg_samples[232] = 16'd968;
ecg_samples[233] = 16'd968;
ecg_samples[234] = 16'd967;
ecg_samples[235] = 16'd969;
ecg_samples[236] = 16'd969;
ecg_samples[237] = 16'd971;
ecg_samples[238] = 16'd970;
ecg_samples[239] = 16'd967;
ecg_samples[240] = 16'd966;
ecg_samples[241] = 16'd968;
ecg_samples[242] = 16'd969;
ecg_samples[243] = 16'd967;
ecg_samples[244] = 16'd968;
ecg_samples[245] = 16'd964;
ecg_samples[246] = 16'd964;
ecg_samples[247] = 16'd963;
ecg_samples[248] = 16'd965;
ecg_samples[249] = 16'd964;
ecg_samples[250] = 16'd962;
ecg_samples[251] = 16'd962;
ecg_samples[252] = 16'd963;
ecg_samples[253] = 16'd965;
ecg_samples[254] = 16'd967;
ecg_samples[255] = 16'd967;
ecg_samples[256] = 16'd966;
ecg_samples[257] = 16'd965;
ecg_samples[258] = 16'd962;
ecg_samples[259] = 16'd966;
ecg_samples[260] = 16'd965;
ecg_samples[261] = 16'd964;
ecg_samples[262] = 16'd963;
ecg_samples[263] = 16'd962;
ecg_samples[264] = 16'd959;
ecg_samples[265] = 16'd962;
ecg_samples[266] = 16'd964;
ecg_samples[267] = 16'd966;
ecg_samples[268] = 16'd962;
ecg_samples[269] = 16'd959;
ecg_samples[270] = 16'd958;
ecg_samples[271] = 16'd961;
ecg_samples[272] = 16'd964;
ecg_samples[273] = 16'd963;
ecg_samples[274] = 16'd962;
ecg_samples[275] = 16'd960;
ecg_samples[276] = 16'd958;
ecg_samples[277] = 16'd959;
ecg_samples[278] = 16'd961;
ecg_samples[279] = 16'd962;
ecg_samples[280] = 16'd963;
ecg_samples[281] = 16'd963;
ecg_samples[282] = 16'd962;
ecg_samples[283] = 16'd964;
ecg_samples[284] = 16'd963;
ecg_samples[285] = 16'd966;
ecg_samples[286] = 16'd964;
ecg_samples[287] = 16'd964;
ecg_samples[288] = 16'd963;
ecg_samples[289] = 16'd963;
ecg_samples[290] = 16'd966;
ecg_samples[291] = 16'd968;
ecg_samples[292] = 16'd965;
ecg_samples[293] = 16'd963;
ecg_samples[294] = 16'd961;
ecg_samples[295] = 16'd963;
ecg_samples[296] = 16'd965;
ecg_samples[297] = 16'd966;
ecg_samples[298] = 16'd968;
ecg_samples[299] = 16'd970;
ecg_samples[300] = 16'd969;
ecg_samples[301] = 16'd969;
ecg_samples[302] = 16'd970;
ecg_samples[303] = 16'd974;
ecg_samples[304] = 16'd974;
ecg_samples[305] = 16'd973;
ecg_samples[306] = 16'd979;
ecg_samples[307] = 16'd980;
ecg_samples[308] = 16'd983;
ecg_samples[309] = 16'd984;
ecg_samples[310] = 16'd983;
ecg_samples[311] = 16'd981;
ecg_samples[312] = 16'd978;
ecg_samples[313] = 16'd980;
ecg_samples[314] = 16'd979;
ecg_samples[315] = 16'd979;
ecg_samples[316] = 16'd979;
ecg_samples[317] = 16'd978;
ecg_samples[318] = 16'd977;
ecg_samples[319] = 16'd976;
ecg_samples[320] = 16'd977;
ecg_samples[321] = 16'd980;
ecg_samples[322] = 16'd982;
ecg_samples[323] = 16'd983;
ecg_samples[324] = 16'd975;
ecg_samples[325] = 16'd967;
ecg_samples[326] = 16'd967;
ecg_samples[327] = 16'd964;
ecg_samples[328] = 16'd962;
ecg_samples[329] = 16'd958;
ecg_samples[330] = 16'd958;
ecg_samples[331] = 16'd959;
ecg_samples[332] = 16'd961;
ecg_samples[333] = 16'd960;
ecg_samples[334] = 16'd961;
ecg_samples[335] = 16'd959;
ecg_samples[336] = 16'd956;
ecg_samples[337] = 16'd955;
ecg_samples[338] = 16'd956;
ecg_samples[339] = 16'd956;
ecg_samples[340] = 16'd954;
ecg_samples[341] = 16'd955;
ecg_samples[342] = 16'd953;
ecg_samples[343] = 16'd958;
ecg_samples[344] = 16'd957;
ecg_samples[345] = 16'd958;
ecg_samples[346] = 16'd960;
ecg_samples[347] = 16'd955;
ecg_samples[348] = 16'd953;
ecg_samples[349] = 16'd956;
ecg_samples[350] = 16'd958;
ecg_samples[351] = 16'd959;
ecg_samples[352] = 16'd958;
ecg_samples[353] = 16'd954;
ecg_samples[354] = 16'd951;
ecg_samples[355] = 16'd952;
ecg_samples[356] = 16'd948;
ecg_samples[357] = 16'd939;
ecg_samples[358] = 16'd935;
ecg_samples[359] = 16'd929;
ecg_samples[360] = 16'd922;
ecg_samples[361] = 16'd917;
ecg_samples[362] = 16'd923;
ecg_samples[363] = 16'd941;
ecg_samples[364] = 16'd964;
ecg_samples[365] = 16'd992;
ecg_samples[366] = 16'd1021;
ecg_samples[367] = 16'd1071;
ecg_samples[368] = 16'd1122;
ecg_samples[369] = 16'd1168;
ecg_samples[370] = 16'd1199;
ecg_samples[371] = 16'd1212;
ecg_samples[372] = 16'd1205;
ecg_samples[373] = 16'd1175;
ecg_samples[374] = 16'd1122;
ecg_samples[375] = 16'd1057;
ecg_samples[376] = 16'd1002;
ecg_samples[377] = 16'd970;
ecg_samples[378] = 16'd946;
ecg_samples[379] = 16'd934;
ecg_samples[380] = 16'd929;
ecg_samples[381] = 16'd933;
ecg_samples[382] = 16'd939;
ecg_samples[383] = 16'd946;
ecg_samples[384] = 16'd946;
ecg_samples[385] = 16'd947;
ecg_samples[386] = 16'd946;
ecg_samples[387] = 16'd948;
ecg_samples[388] = 16'd948;
ecg_samples[389] = 16'd948;
ecg_samples[390] = 16'd945;
ecg_samples[391] = 16'd947;
ecg_samples[392] = 16'd947;
ecg_samples[393] = 16'd947;
ecg_samples[394] = 16'd949;
ecg_samples[395] = 16'd945;
ecg_samples[396] = 16'd942;
ecg_samples[397] = 16'd942;
ecg_samples[398] = 16'd944;
ecg_samples[399] = 16'd945;
ecg_samples[400] = 16'd946;
ecg_samples[401] = 16'd943;
ecg_samples[402] = 16'd945;
ecg_samples[403] = 16'd947;
ecg_samples[404] = 16'd949;
ecg_samples[405] = 16'd946;
ecg_samples[406] = 16'd946;
ecg_samples[407] = 16'd943;
ecg_samples[408] = 16'd942;
ecg_samples[409] = 16'd942;
ecg_samples[410] = 16'd946;
ecg_samples[411] = 16'd946;
ecg_samples[412] = 16'd945;
ecg_samples[413] = 16'd943;
ecg_samples[414] = 16'd941;
ecg_samples[415] = 16'd944;
ecg_samples[416] = 16'd942;
ecg_samples[417] = 16'd943;
ecg_samples[418] = 16'd942;
ecg_samples[419] = 16'd941;
ecg_samples[420] = 16'd942;
ecg_samples[421] = 16'd944;
ecg_samples[422] = 16'd944;
ecg_samples[423] = 16'd945;
ecg_samples[424] = 16'd946;
ecg_samples[425] = 16'd943;
ecg_samples[426] = 16'd942;
ecg_samples[427] = 16'd946;
ecg_samples[428] = 16'd946;
ecg_samples[429] = 16'd947;
ecg_samples[430] = 16'd947;
ecg_samples[431] = 16'd942;
ecg_samples[432] = 16'd943;
ecg_samples[433] = 16'd945;
ecg_samples[434] = 16'd946;
ecg_samples[435] = 16'd949;
ecg_samples[436] = 16'd946;
ecg_samples[437] = 16'd945;
ecg_samples[438] = 16'd942;
ecg_samples[439] = 16'd944;
ecg_samples[440] = 16'd946;
ecg_samples[441] = 16'd946;
ecg_samples[442] = 16'd947;
ecg_samples[443] = 16'd943;
ecg_samples[444] = 16'd941;
ecg_samples[445] = 16'd941;
ecg_samples[446] = 16'd944;
ecg_samples[447] = 16'd945;
ecg_samples[448] = 16'd943;
ecg_samples[449] = 16'd941;
ecg_samples[450] = 16'd940;
ecg_samples[451] = 16'd940;
ecg_samples[452] = 16'd942;
ecg_samples[453] = 16'd941;
ecg_samples[454] = 16'd939;
ecg_samples[455] = 16'd940;
ecg_samples[456] = 16'd937;
ecg_samples[457] = 16'd938;
ecg_samples[458] = 16'd938;
ecg_samples[459] = 16'd940;
ecg_samples[460] = 16'd938;
ecg_samples[461] = 16'd934;
ecg_samples[462] = 16'd933;
ecg_samples[463] = 16'd934;
ecg_samples[464] = 16'd937;
ecg_samples[465] = 16'd935;
ecg_samples[466] = 16'd934;
ecg_samples[467] = 16'd933;
ecg_samples[468] = 16'd930;
ecg_samples[469] = 16'd932;
ecg_samples[470] = 16'd933;
ecg_samples[471] = 16'd934;
ecg_samples[472] = 16'd933;
ecg_samples[473] = 16'd930;
ecg_samples[474] = 16'd929;
ecg_samples[475] = 16'd932;
ecg_samples[476] = 16'd934;
ecg_samples[477] = 16'd935;
ecg_samples[478] = 16'd936;
ecg_samples[479] = 16'd937;
ecg_samples[480] = 16'd936;
ecg_samples[481] = 16'd942;
ecg_samples[482] = 16'd945;
ecg_samples[483] = 16'd950;
ecg_samples[484] = 16'd951;
ecg_samples[485] = 16'd952;
ecg_samples[486] = 16'd951;
ecg_samples[487] = 16'd956;
ecg_samples[488] = 16'd959;
ecg_samples[489] = 16'd961;
ecg_samples[490] = 16'd960;
ecg_samples[491] = 16'd958;
ecg_samples[492] = 16'd958;
ecg_samples[493] = 16'd960;
ecg_samples[494] = 16'd962;
ecg_samples[495] = 16'd964;
ecg_samples[496] = 16'd964;
ecg_samples[497] = 16'd960;
ecg_samples[498] = 16'd960;
ecg_samples[499] = 16'd961;
ecg_samples[500] = 16'd963;
ecg_samples[501] = 16'd963;
ecg_samples[502] = 16'd965;
ecg_samples[503] = 16'd960;
ecg_samples[504] = 16'd958;
ecg_samples[505] = 16'd963;
ecg_samples[506] = 16'd962;
ecg_samples[507] = 16'd964;
ecg_samples[508] = 16'd964;
ecg_samples[509] = 16'd960;
ecg_samples[510] = 16'd959;
ecg_samples[511] = 16'd962;
ecg_samples[512] = 16'd963;
ecg_samples[513] = 16'd961;
ecg_samples[514] = 16'd963;
ecg_samples[515] = 16'd961;
ecg_samples[516] = 16'd961;
ecg_samples[517] = 16'd962;
ecg_samples[518] = 16'd965;
ecg_samples[519] = 16'd966;
ecg_samples[520] = 16'd963;
ecg_samples[521] = 16'd962;
ecg_samples[522] = 16'd960;
ecg_samples[523] = 16'd961;
ecg_samples[524] = 16'd964;
ecg_samples[525] = 16'd961;
ecg_samples[526] = 16'd961;
ecg_samples[527] = 16'd961;
ecg_samples[528] = 16'd958;
ecg_samples[529] = 16'd961;
ecg_samples[530] = 16'd960;
ecg_samples[531] = 16'd961;
ecg_samples[532] = 16'd959;
ecg_samples[533] = 16'd957;
ecg_samples[534] = 16'd956;
ecg_samples[535] = 16'd957;
ecg_samples[536] = 16'd957;
ecg_samples[537] = 16'd958;
ecg_samples[538] = 16'd959;
ecg_samples[539] = 16'd955;
ecg_samples[540] = 16'd954;
ecg_samples[541] = 16'd955;
ecg_samples[542] = 16'd957;
ecg_samples[543] = 16'd958;
ecg_samples[544] = 16'd958;
ecg_samples[545] = 16'd955;
ecg_samples[546] = 16'd955;
ecg_samples[547] = 16'd955;
ecg_samples[548] = 16'd960;
ecg_samples[549] = 16'd958;
ecg_samples[550] = 16'd957;
ecg_samples[551] = 16'd956;
ecg_samples[552] = 16'd953;
ecg_samples[553] = 16'd957;
ecg_samples[554] = 16'd958;
ecg_samples[555] = 16'd958;
ecg_samples[556] = 16'd957;
ecg_samples[557] = 16'd953;
ecg_samples[558] = 16'd952;
ecg_samples[559] = 16'd953;
ecg_samples[560] = 16'd954;
ecg_samples[561] = 16'd956;
ecg_samples[562] = 16'd955;
ecg_samples[563] = 16'd955;
ecg_samples[564] = 16'd955;
ecg_samples[565] = 16'd955;
ecg_samples[566] = 16'd958;
ecg_samples[567] = 16'd958;
ecg_samples[568] = 16'd957;
ecg_samples[569] = 16'd955;
ecg_samples[570] = 16'd954;
ecg_samples[571] = 16'd954;
ecg_samples[572] = 16'd956;
ecg_samples[573] = 16'd958;
ecg_samples[574] = 16'd955;
ecg_samples[575] = 16'd955;
ecg_samples[576] = 16'd953;
ecg_samples[577] = 16'd954;
ecg_samples[578] = 16'd956;
ecg_samples[579] = 16'd958;
ecg_samples[580] = 16'd956;
ecg_samples[581] = 16'd956;
ecg_samples[582] = 16'd956;
ecg_samples[583] = 16'd958;
ecg_samples[584] = 16'd957;
ecg_samples[585] = 16'd958;
ecg_samples[586] = 16'd957;
ecg_samples[587] = 16'd955;
ecg_samples[588] = 16'd955;
ecg_samples[589] = 16'd956;
ecg_samples[590] = 16'd958;
ecg_samples[591] = 16'd961;
ecg_samples[592] = 16'd965;
ecg_samples[593] = 16'd964;
ecg_samples[594] = 16'd965;
ecg_samples[595] = 16'd967;
ecg_samples[596] = 16'd969;
ecg_samples[597] = 16'd971;
ecg_samples[598] = 16'd971;
ecg_samples[599] = 16'd971;
ecg_samples[600] = 16'd973;
ecg_samples[601] = 16'd974;
ecg_samples[602] = 16'd976;
ecg_samples[603] = 16'd979;
ecg_samples[604] = 16'd981;
ecg_samples[605] = 16'd976;
ecg_samples[606] = 16'd975;
ecg_samples[607] = 16'd976;
ecg_samples[608] = 16'd975;
ecg_samples[609] = 16'd977;
ecg_samples[610] = 16'd975;
ecg_samples[611] = 16'd974;
ecg_samples[612] = 16'd969;
ecg_samples[613] = 16'd969;
ecg_samples[614] = 16'd971;
ecg_samples[615] = 16'd974;
ecg_samples[616] = 16'd979;
ecg_samples[617] = 16'd980;
ecg_samples[618] = 16'd978;
ecg_samples[619] = 16'd971;
ecg_samples[620] = 16'd970;
ecg_samples[621] = 16'd968;
ecg_samples[622] = 16'd967;
ecg_samples[623] = 16'd963;
ecg_samples[624] = 16'd960;
ecg_samples[625] = 16'd956;
ecg_samples[626] = 16'd958;
ecg_samples[627] = 16'd957;
ecg_samples[628] = 16'd957;
ecg_samples[629] = 16'd953;
ecg_samples[630] = 16'd950;
ecg_samples[631] = 16'd952;
ecg_samples[632] = 16'd955;
ecg_samples[633] = 16'd954;
ecg_samples[634] = 16'd953;
ecg_samples[635] = 16'd951;
ecg_samples[636] = 16'd949;
ecg_samples[637] = 16'd948;
ecg_samples[638] = 16'd950;
ecg_samples[639] = 16'd951;
ecg_samples[640] = 16'd951;
ecg_samples[641] = 16'd948;
ecg_samples[642] = 16'd947;
ecg_samples[643] = 16'd948;
ecg_samples[644] = 16'd949;
ecg_samples[645] = 16'd953;
ecg_samples[646] = 16'd950;
ecg_samples[647] = 16'd946;
ecg_samples[648] = 16'd943;
ecg_samples[649] = 16'd942;
ecg_samples[650] = 16'd937;
ecg_samples[651] = 16'd931;
ecg_samples[652] = 16'd926;
ecg_samples[653] = 16'd920;
ecg_samples[654] = 16'd913;
ecg_samples[655] = 16'd910;
ecg_samples[656] = 16'd919;
ecg_samples[657] = 16'd943;
ecg_samples[658] = 16'd974;
ecg_samples[659] = 16'd1006;
ecg_samples[660] = 16'd1048;
ecg_samples[661] = 16'd1106;
ecg_samples[662] = 16'd1162;
ecg_samples[663] = 16'd1201;
ecg_samples[664] = 16'd1216;
ecg_samples[665] = 16'd1194;
ecg_samples[666] = 16'd1128;
ecg_samples[667] = 16'd1034;
ecg_samples[668] = 16'd960;
ecg_samples[669] = 16'd924;
ecg_samples[670] = 16'd923;
ecg_samples[671] = 16'd935;
ecg_samples[672] = 16'd941;
ecg_samples[673] = 16'd945;
ecg_samples[674] = 16'd946;
ecg_samples[675] = 16'd945;
ecg_samples[676] = 16'd946;
ecg_samples[677] = 16'd945;
ecg_samples[678] = 16'd943;
ecg_samples[679] = 16'd945;
ecg_samples[680] = 16'd943;
ecg_samples[681] = 16'd946;
ecg_samples[682] = 16'd945;
ecg_samples[683] = 16'd945;
ecg_samples[684] = 16'd942;
ecg_samples[685] = 16'd943;
ecg_samples[686] = 16'd944;
ecg_samples[687] = 16'd944;
ecg_samples[688] = 16'd941;
ecg_samples[689] = 16'd943;
ecg_samples[690] = 16'd940;
ecg_samples[691] = 16'd941;
ecg_samples[692] = 16'd943;
ecg_samples[693] = 16'd943;
ecg_samples[694] = 16'd940;
ecg_samples[695] = 16'd940;
ecg_samples[696] = 16'd937;
ecg_samples[697] = 16'd940;
ecg_samples[698] = 16'd942;
ecg_samples[699] = 16'd942;
ecg_samples[700] = 16'd943;
ecg_samples[701] = 16'd939;
ecg_samples[702] = 16'd938;
ecg_samples[703] = 16'd940;
ecg_samples[704] = 16'd941;
ecg_samples[705] = 16'd942;
ecg_samples[706] = 16'd942;
ecg_samples[707] = 16'd939;
ecg_samples[708] = 16'd940;
ecg_samples[709] = 16'd944;
ecg_samples[710] = 16'd945;
ecg_samples[711] = 16'd944;
ecg_samples[712] = 16'd944;
ecg_samples[713] = 16'd945;
ecg_samples[714] = 16'd941;
ecg_samples[715] = 16'd943;
ecg_samples[716] = 16'd946;
ecg_samples[717] = 16'd944;
ecg_samples[718] = 16'd944;
ecg_samples[719] = 16'd941;
ecg_samples[720] = 16'd939;
ecg_samples[721] = 16'd939;
ecg_samples[722] = 16'd941;
ecg_samples[723] = 16'd941;
ecg_samples[724] = 16'd942;
ecg_samples[725] = 16'd939;
ecg_samples[726] = 16'd939;
ecg_samples[727] = 16'd940;
ecg_samples[728] = 16'd941;
ecg_samples[729] = 16'd944;
ecg_samples[730] = 16'd944;
ecg_samples[731] = 16'd942;
ecg_samples[732] = 16'd939;
ecg_samples[733] = 16'd942;
ecg_samples[734] = 16'd943;
ecg_samples[735] = 16'd945;
ecg_samples[736] = 16'd944;
ecg_samples[737] = 16'd944;
ecg_samples[738] = 16'd943;
ecg_samples[739] = 16'd947;
ecg_samples[740] = 16'd944;
ecg_samples[741] = 16'd946;
ecg_samples[742] = 16'd946;
ecg_samples[743] = 16'd944;
ecg_samples[744] = 16'd941;
ecg_samples[745] = 16'd943;
ecg_samples[746] = 16'd943;
ecg_samples[747] = 16'd942;
ecg_samples[748] = 16'd941;
ecg_samples[749] = 16'd940;
ecg_samples[750] = 16'd940;
ecg_samples[751] = 16'd939;
ecg_samples[752] = 16'd941;
ecg_samples[753] = 16'd941;
ecg_samples[754] = 16'd942;
ecg_samples[755] = 16'd937;
ecg_samples[756] = 16'd938;
ecg_samples[757] = 16'd937;
ecg_samples[758] = 16'd940;
ecg_samples[759] = 16'd940;
ecg_samples[760] = 16'd940;
ecg_samples[761] = 16'd940;
ecg_samples[762] = 16'd939;
ecg_samples[763] = 16'd939;
ecg_samples[764] = 16'd941;
ecg_samples[765] = 16'd945;
ecg_samples[766] = 16'd945;
ecg_samples[767] = 16'd946;
ecg_samples[768] = 16'd949;
ecg_samples[769] = 16'd952;
ecg_samples[770] = 16'd956;
ecg_samples[771] = 16'd957;
ecg_samples[772] = 16'd958;
ecg_samples[773] = 16'd957;
ecg_samples[774] = 16'd957;
ecg_samples[775] = 16'd959;
ecg_samples[776] = 16'd960;
ecg_samples[777] = 16'd963;
ecg_samples[778] = 16'd963;
ecg_samples[779] = 16'd961;
ecg_samples[780] = 16'd962;
ecg_samples[781] = 16'd963;
ecg_samples[782] = 16'd964;
ecg_samples[783] = 16'd964;
ecg_samples[784] = 16'd964;
ecg_samples[785] = 16'd962;
ecg_samples[786] = 16'd962;
ecg_samples[787] = 16'd962;
ecg_samples[788] = 16'd961;
ecg_samples[789] = 16'd964;
ecg_samples[790] = 16'd963;
ecg_samples[791] = 16'd961;
ecg_samples[792] = 16'd960;
ecg_samples[793] = 16'd959;
ecg_samples[794] = 16'd962;
ecg_samples[795] = 16'd963;
ecg_samples[796] = 16'd963;
ecg_samples[797] = 16'd960;
ecg_samples[798] = 16'd959;
ecg_samples[799] = 16'd963;
ecg_samples[800] = 16'd962;
ecg_samples[801] = 16'd965;
ecg_samples[802] = 16'd962;
ecg_samples[803] = 16'd959;
ecg_samples[804] = 16'd958;
ecg_samples[805] = 16'd960;
ecg_samples[806] = 16'd960;
ecg_samples[807] = 16'd960;
ecg_samples[808] = 16'd959;
ecg_samples[809] = 16'd954;
ecg_samples[810] = 16'd954;
ecg_samples[811] = 16'd956;
ecg_samples[812] = 16'd957;
ecg_samples[813] = 16'd958;
ecg_samples[814] = 16'd957;
ecg_samples[815] = 16'd956;
ecg_samples[816] = 16'd952;
ecg_samples[817] = 16'd954;
ecg_samples[818] = 16'd954;
ecg_samples[819] = 16'd953;
ecg_samples[820] = 16'd952;
ecg_samples[821] = 16'd953;
ecg_samples[822] = 16'd951;
ecg_samples[823] = 16'd953;
ecg_samples[824] = 16'd954;
ecg_samples[825] = 16'd956;
ecg_samples[826] = 16'd953;
ecg_samples[827] = 16'd954;
ecg_samples[828] = 16'd951;
ecg_samples[829] = 16'd951;
ecg_samples[830] = 16'd954;
ecg_samples[831] = 16'd953;
ecg_samples[832] = 16'd954;
ecg_samples[833] = 16'd950;
ecg_samples[834] = 16'd948;
ecg_samples[835] = 16'd950;
ecg_samples[836] = 16'd952;
ecg_samples[837] = 16'd951;
ecg_samples[838] = 16'd952;
ecg_samples[839] = 16'd951;
ecg_samples[840] = 16'd948;
ecg_samples[841] = 16'd950;
ecg_samples[842] = 16'd951;
ecg_samples[843] = 16'd954;
ecg_samples[844] = 16'd954;
ecg_samples[845] = 16'd954;
ecg_samples[846] = 16'd950;
ecg_samples[847] = 16'd951;
ecg_samples[848] = 16'd955;
ecg_samples[849] = 16'd955;
ecg_samples[850] = 16'd956;
ecg_samples[851] = 16'd953;
ecg_samples[852] = 16'd951;
ecg_samples[853] = 16'd952;
ecg_samples[854] = 16'd953;
ecg_samples[855] = 16'd953;
ecg_samples[856] = 16'd953;
ecg_samples[857] = 16'd949;
ecg_samples[858] = 16'd947;
ecg_samples[859] = 16'd953;
ecg_samples[860] = 16'd952;
ecg_samples[861] = 16'd953;
ecg_samples[862] = 16'd952;
ecg_samples[863] = 16'd952;
ecg_samples[864] = 16'd950;
ecg_samples[865] = 16'd952;
ecg_samples[866] = 16'd955;
ecg_samples[867] = 16'd953;
ecg_samples[868] = 16'd955;
ecg_samples[869] = 16'd955;
ecg_samples[870] = 16'd955;
ecg_samples[871] = 16'd956;
ecg_samples[872] = 16'd962;
ecg_samples[873] = 16'd963;
ecg_samples[874] = 16'd963;
ecg_samples[875] = 16'd962;
ecg_samples[876] = 16'd963;
ecg_samples[877] = 16'd966;
ecg_samples[878] = 16'd967;
ecg_samples[879] = 16'd969;
ecg_samples[880] = 16'd968;
ecg_samples[881] = 16'd968;
ecg_samples[882] = 16'd969;
ecg_samples[883] = 16'd971;
ecg_samples[884] = 16'd973;
ecg_samples[885] = 16'd975;
ecg_samples[886] = 16'd972;
ecg_samples[887] = 16'd971;
ecg_samples[888] = 16'd969;
ecg_samples[889] = 16'd968;
ecg_samples[890] = 16'd971;
ecg_samples[891] = 16'd970;
ecg_samples[892] = 16'd969;
ecg_samples[893] = 16'd968;
ecg_samples[894] = 16'd969;
ecg_samples[895] = 16'd968;
ecg_samples[896] = 16'd969;
ecg_samples[897] = 16'd971;
ecg_samples[898] = 16'd973;
ecg_samples[899] = 16'd976;
ecg_samples[900] = 16'd972;
ecg_samples[901] = 16'd968;
ecg_samples[902] = 16'd962;
ecg_samples[903] = 16'd962;
ecg_samples[904] = 16'd955;
ecg_samples[905] = 16'd952;
ecg_samples[906] = 16'd948;
ecg_samples[907] = 16'd947;
ecg_samples[908] = 16'd948;
ecg_samples[909] = 16'd950;
ecg_samples[910] = 16'd949;
ecg_samples[911] = 16'd947;
ecg_samples[912] = 16'd946;
ecg_samples[913] = 16'd945;
ecg_samples[914] = 16'd947;
ecg_samples[915] = 16'd947;
ecg_samples[916] = 16'd947;
ecg_samples[917] = 16'd945;
ecg_samples[918] = 16'd943;
ecg_samples[919] = 16'd944;
ecg_samples[920] = 16'd949;
ecg_samples[921] = 16'd949;
ecg_samples[922] = 16'd946;
ecg_samples[923] = 16'd945;
ecg_samples[924] = 16'd941;
ecg_samples[925] = 16'd943;
ecg_samples[926] = 16'd944;
ecg_samples[927] = 16'd946;
ecg_samples[928] = 16'd943;
ecg_samples[929] = 16'd939;
ecg_samples[930] = 16'd932;
ecg_samples[931] = 16'd929;
ecg_samples[932] = 16'd923;
ecg_samples[933] = 16'd922;
ecg_samples[934] = 16'd919;
ecg_samples[935] = 16'd916;
ecg_samples[936] = 16'd904;
ecg_samples[937] = 16'd895;
ecg_samples[938] = 16'd898;
ecg_samples[939] = 16'd909;
ecg_samples[940] = 16'd925;
ecg_samples[941] = 16'd947;
ecg_samples[942] = 16'd970;
ecg_samples[943] = 16'd1001;
ecg_samples[944] = 16'd1042;
ecg_samples[945] = 16'd1098;
ecg_samples[946] = 16'd1151;
ecg_samples[947] = 16'd1186;
ecg_samples[948] = 16'd1196;
ecg_samples[949] = 16'd1178;
ecg_samples[950] = 16'd1119;
ecg_samples[951] = 16'd1037;
ecg_samples[952] = 16'd963;
ecg_samples[953] = 16'd924;
ecg_samples[954] = 16'd920;
ecg_samples[955] = 16'd929;
ecg_samples[956] = 16'd942;
ecg_samples[957] = 16'd946;
ecg_samples[958] = 16'd946;
ecg_samples[959] = 16'd944;
ecg_samples[960] = 16'd942;
ecg_samples[961] = 16'd943;
ecg_samples[962] = 16'd947;
ecg_samples[963] = 16'd946;
ecg_samples[964] = 16'd945;
ecg_samples[965] = 16'd943;
ecg_samples[966] = 16'd942;
ecg_samples[967] = 16'd943;
ecg_samples[968] = 16'd944;
ecg_samples[969] = 16'd946;
ecg_samples[970] = 16'd945;
ecg_samples[971] = 16'd942;
ecg_samples[972] = 16'd941;
ecg_samples[973] = 16'd942;
ecg_samples[974] = 16'd945;
ecg_samples[975] = 16'd943;
ecg_samples[976] = 16'd942;
ecg_samples[977] = 16'd943;
ecg_samples[978] = 16'd943;
ecg_samples[979] = 16'd942;
ecg_samples[980] = 16'd946;
ecg_samples[981] = 16'd947;
ecg_samples[982] = 16'd946;
ecg_samples[983] = 16'd945;
ecg_samples[984] = 16'd944;
ecg_samples[985] = 16'd944;
ecg_samples[986] = 16'd944;
ecg_samples[987] = 16'd945;
ecg_samples[988] = 16'd945;
ecg_samples[989] = 16'd943;
ecg_samples[990] = 16'd943;
ecg_samples[991] = 16'd944;
ecg_samples[992] = 16'd945;
ecg_samples[993] = 16'd947;
ecg_samples[994] = 16'd949;
ecg_samples[995] = 16'd947;
ecg_samples[996] = 16'd945;
ecg_samples[997] = 16'd946;
ecg_samples[998] = 16'd947;
ecg_samples[999] = 16'd949;

// Add powerline interference and baseline wander
for (i = 0; i < 1000; i=i+1) begin
  ecg_samples[i] = ecg_samples[i] + 16'd2 * $sin(2 * 3.14159 * 50 * i / 1000); // add 50Hz powerline interference
  ecg_samples[i] = ecg_samples[i] + 16'd5 * $sin(2 * 3.14159 * 0.5 * i / 1000); // add baseline wander
end

clk = 0;
reset = 1;
sample = 0;
#100;
reset = 0;

for (i = 0; i < 1000; i=i+1) begin
sample = ecg_samples[i];
#10;
clk = 1;
#10;
clk = 0;
$display(" %d", result);
end
end
endmodule

